// `include "VAPE_immutability.v"
// `include "VAPE_atomicity.v"
// `include "VAPE_output_protection.v"
// `include "VAPE_EXEC_flag.v"
// `include "VAPE_boundary.v"
// `include "VAPE_reset.v"
// `include "VAPE_irq_dma.v"

`include "log_monitor.v"
`include "slice_monitor.v"
`include "branch_monitor.v"
`include "boundary_monitor.v"
`include "loop_monitor.v"
`include "logger.v"

`ifdef OMSP_NO_INCLUDE
`else
`include "openMSP430_defines.v"
`endif

module cflow (
    clk,
    pc,
    pc_nxt,
    
    data_wr,
    data_addr,
    
    dma_addr,
    dma_en,
    
    puc,

    ER_min,
    ER_max,

    irq_ta0,
    irq,
    gie,
    
    e_state,
    inst_so,
    inst_type,
    inst_ad,
    inst_as,
    inst_jmp,
    
    cflow_hw_wen,
    cflow_log_ptr,
    cflow_src,
    cflow_dest,
    
    reset,
    flush_log,
    boot,
    ER_done,

    flush_slice,
    top_slice,
    bottom_slice
);
input           clk;
input   [15:0]  pc;
input   [15:0]  pc_nxt;
input           data_wr;
input   [15:0]  data_addr;
input   [15:0]  dma_addr;
input           dma_en;
input   [15:0]  ER_min;
input   [15:0]  ER_max;
input           puc;
input           irq_ta0;
input           irq;
input           gie;
input   [3:0]   e_state;
input   [7:0]   inst_so;
input   [2:0]   inst_type;
input   [7:0]   inst_ad;
input   [7:0]   inst_as;
input   [7:0]   inst_jmp;
// 
output          cflow_hw_wen;
output  [15:0]  cflow_log_ptr;
output  [15:0]  cflow_src;
output  [15:0]  cflow_dest; 
output          reset;
output          flush_log;
output          boot;
output          ER_done;
// outputs from slice monitor
output          flush_slice;
output  [15:0]  top_slice;
output  [15:0]  bottom_slice; 




//// log size in WORDS\
parameter LOG_SIZE = `LOG_SIZE/2;

// parameter LOG_SIZE = 16'h0080; // 256
// parameter LOG_SIZE = 16'h0100; // 512
//parameter LOG_SIZE = 16'h0200; // 1024
// parameter LOG_SIZE = 16'h0400; // 2048
//parameter LOG_SIZE = 16'h0800;   // total words for 4096 bytes cflog  (4kb)
//parameter LOG_SIZE = 16'h1000;   // total words for 8192 bytes cflog  (8kb)
//parameter LOG_SIZE = 16'h1800;   // total words for 12288 bytes cflog  (12kb)
//
parameter TCB_max = 16'hdffe; 
parameter RESET_addr = 16'he000;
parameter PMEM_min = 16'he03e;

reg tcb_boot_done = 0;
reg [15:0] prev_pc;
// wire [15:0] cflow_log_prev_ptr;
wire [31:0] loop_ctr;
wire loop_detect_out;
wire pc_in_ER = (pc >= ER_min) && (pc <= ER_max) && (ER_min != 0) && (ER_max != 0);
wire caramel_timer = irq_ta0 & pc_in_ER;
wire acfa_nmi = caramel_timer | flush_log | flush_slice | ER_done | boot;
// wire pc_TCB_exit = (pc == TCB_max);

// boundary_monitor #(
//     .LOG_SIZE (LOG_SIZE)) 
// boundary_monitor_0 ( // Boundary Protection
//     .clk        (clk),
//     .pc         (pc),
//     .data_addr  (data_addr),
//     .data_en    (data_wr),
//     .dma_addr   (dma_addr),
//     .dma_en     (dma_en),
//     .ER_min     (ER_min),
//     .ER_max     (ER_max),
//     .reset      (reset) 
// );

log_monitor #(
    .LOG_SIZE (LOG_SIZE)
) 
log_monitor_0 (
    .clk        (clk),
    .pc         (pc),
    .pc_nxt     (pc_nxt),    
    .ER_min     (ER_min),
    .ER_max     (ER_max),
    .irq        (irq),
    .reset      (puc),
    .loop_detect    (loop_detect_out),
    .branch_detect  (branch_detect),
    .top_slice      (top_slice),

    // outputs
    .flush      (flush_log),
    .hw_wr_en       (cflow_hw_wen),
    .cflow_log_ptr  (cflow_log_ptr)
);

branch_monitor #(
    .LOG_SIZE (LOG_SIZE)
)
branch_monitor_0( //Branch Monitor
    
    .clk            (clk),    
    .pc             (pc),     
    .ER_min         (ER_min),
    .ER_max         (ER_max),
    .acfa_nmi   (acfa_nmi),
    .irq        (irq),
    .gie        (gie),

    .e_state    (e_state),
    .inst_so    (inst_so),
    .inst_type  (inst_type),
    .inst_ad    (inst_ad),
    .inst_as    (inst_as),
    .inst_jmp   (inst_jmp),
    
    .branch_detect (branch_detect)
);


slice_monitor #(
    .LOG_SIZE (LOG_SIZE)
) 
slice_monitor_0 (
    .clk           (clk),
    .pc            (pc),
    .pc_nxt        (pc_nxt),
    
    .ER_done       (ER_done),
    .ER_min        (ER_min),
    .ER_max        (ER_max),
 
    .irq           (irq),
    .reset         (puc),
    .cflow_log_ptr (cflow_log_ptr),

    .flush          (flush_slice),
    .top_slice      (top_slice),
    .bottom_slice   (bottom_slice)
);

always @(posedge clk)
begin
    prev_pc <= pc;  
end

loop_monitor loop_monitor_0(
    .clk            (clk),    
    .pc             (pc),
    .pc_nxt         (pc_nxt),
    // .prev_pc        (prev_pc),
    
    // .acfa_nmi       (acfa_nmi),
    // .hw_wr_en       (cflow_hw_wen),
    .branch_detect  (branch_detect),
    
    .loop_detect    (loop_detect_out),
    .loop_ctr       (loop_ctr)
);

logger logger_0(
    // .clk            (clk),
    .pc             (pc),
    .prev_pc        (prev_pc),
    
    .loop_detect    (loop_detect_out),
    .loop_ctr       (loop_ctr),
    .cflow_src      (cflow_src),
    .cflow_dest     (cflow_dest)
);

always @(posedge clk) 
begin
   if(pc == TCB_max)
      tcb_boot_done <= 1'b1;
   else if(reset)
      tcb_boot_done <= 1'b0;
   else
      tcb_boot_done <= tcb_boot_done;
end

assign ER_done = (pc == ER_max) & tcb_boot_done;
assign boot = (pc == PMEM_min);

endmodule //cflow
